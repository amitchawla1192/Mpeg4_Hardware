-- VHDL global package produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
package ahir_system_global_package is -- 
  constant job_base_address : std_logic_vector(7 downto 0) := "00000000";
  constant mempool_base_address : std_logic_vector(0 downto 0) := "0";
  -- 
end package ahir_system_global_package;
